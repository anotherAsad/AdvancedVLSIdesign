// serves to load the coefficients for synthesis.
module coeff_broadcaster;
	reg  [15:0] fir_coeff [0:`FILTER_SIZE-1];

		initial begin
		fir_coeff[0] = 16'h0;
		fir_coeff[1] = 16'hFFFF;
		fir_coeff[2] = 16'hFFFE;
		fir_coeff[3] = 16'hFFFB;
		fir_coeff[4] = 16'hFFF8;
		fir_coeff[5] = 16'hFFF4;
		fir_coeff[6] = 16'hFFF2;
		fir_coeff[7] = 16'hFFF1;
		fir_coeff[8] = 16'hFFF2;
		fir_coeff[9] = 16'hFFF6;
		fir_coeff[10] = 16'hFFFC;
		fir_coeff[11] = 16'h2;
		fir_coeff[12] = 16'h7;
		fir_coeff[13] = 16'h9;
		fir_coeff[14] = 16'h8;
		fir_coeff[15] = 16'h4;
		fir_coeff[16] = 16'hFFFE;
		fir_coeff[17] = 16'hFFF9;
		fir_coeff[18] = 16'hFFF7;
		fir_coeff[19] = 16'hFFF8;
		fir_coeff[20] = 16'hFFFD;
		fir_coeff[21] = 16'h3;
		fir_coeff[22] = 16'h9;
		fir_coeff[23] = 16'hB;
		fir_coeff[24] = 16'h8;
		fir_coeff[25] = 16'h2;
		fir_coeff[26] = 16'hFFFB;
		fir_coeff[27] = 16'hFFF5;
		fir_coeff[28] = 16'hFFF3;
		fir_coeff[29] = 16'hFFF7;
		fir_coeff[30] = 16'hFFFF;
		fir_coeff[31] = 16'h8;
		fir_coeff[32] = 16'hE;
		fir_coeff[33] = 16'hF;
		fir_coeff[34] = 16'h9;
		fir_coeff[35] = 16'hFFFF;
		fir_coeff[36] = 16'hFFF4;
		fir_coeff[37] = 16'hFFEE;
		fir_coeff[38] = 16'hFFEF;
		fir_coeff[39] = 16'hFFF8;
		fir_coeff[40] = 16'h5;
		fir_coeff[41] = 16'h11;
		fir_coeff[42] = 16'h17;
		fir_coeff[43] = 16'h13;
		fir_coeff[44] = 16'h7;
		fir_coeff[45] = 16'hFFF7;
		fir_coeff[46] = 16'hFFE9;
		fir_coeff[47] = 16'hFFE5;
		fir_coeff[48] = 16'hFFEB;
		fir_coeff[49] = 16'hFFFC;
		fir_coeff[50] = 16'hF;
		fir_coeff[51] = 16'h1E;
		fir_coeff[52] = 16'h20;
		fir_coeff[53] = 16'h15;
		fir_coeff[54] = 16'h0;
		fir_coeff[55] = 16'hFFE9;
		fir_coeff[56] = 16'hFFDA;
		fir_coeff[57] = 16'hFFDB;
		fir_coeff[58] = 16'hFFEC;
		fir_coeff[59] = 16'h7;
		fir_coeff[60] = 16'h22;
		fir_coeff[61] = 16'h30;
		fir_coeff[62] = 16'h2A;
		fir_coeff[63] = 16'h11;
		fir_coeff[64] = 16'hFFEF;
		fir_coeff[65] = 16'hFFD1;
		fir_coeff[66] = 16'hFFC6;
		fir_coeff[67] = 16'hFFD3;
		fir_coeff[68] = 16'hFFF5;
		fir_coeff[69] = 16'h1F;
		fir_coeff[70] = 16'h3F;
		fir_coeff[71] = 16'h46;
		fir_coeff[72] = 16'h2F;
		fir_coeff[73] = 16'h1;
		fir_coeff[74] = 16'hFFCE;
		fir_coeff[75] = 16'hFFAC;
		fir_coeff[76] = 16'hFFAC;
		fir_coeff[77] = 16'hFFD2;
		fir_coeff[78] = 16'h10;
		fir_coeff[79] = 16'h4D;
		fir_coeff[80] = 16'h6F;
		fir_coeff[81] = 16'h63;
		fir_coeff[82] = 16'h2A;
		fir_coeff[83] = 16'hFFD6;
		fir_coeff[84] = 16'hFF8B;
		fir_coeff[85] = 16'hFF6A;
		fir_coeff[86] = 16'hFF88;
		fir_coeff[87] = 16'hFFE2;
		fir_coeff[88] = 16'h58;
		fir_coeff[89] = 16'hB9;
		fir_coeff[90] = 16'hD7;
		fir_coeff[91] = 16'h97;
		fir_coeff[92] = 16'h2;
		fir_coeff[93] = 16'hFF47;
		fir_coeff[94] = 16'hFEB3;
		fir_coeff[95] = 16'hFE93;
		fir_coeff[96] = 16'hFF1E;
		fir_coeff[97] = 16'h5D;
		fir_coeff[98] = 16'h222;
		fir_coeff[99] = 16'h40E;
		fir_coeff[100] = 16'h5B0;
		fir_coeff[101] = 16'h69F;
		fir_coeff[102] = 16'h69F;
		fir_coeff[103] = 16'h5B0;
		fir_coeff[104] = 16'h40E;
		fir_coeff[105] = 16'h222;
		fir_coeff[106] = 16'h5D;
		fir_coeff[107] = 16'hFF1E;
		fir_coeff[108] = 16'hFE93;
		fir_coeff[109] = 16'hFEB3;
		fir_coeff[110] = 16'hFF47;
		fir_coeff[111] = 16'h2;
		fir_coeff[112] = 16'h97;
		fir_coeff[113] = 16'hD7;
		fir_coeff[114] = 16'hB9;
		fir_coeff[115] = 16'h58;
		fir_coeff[116] = 16'hFFE2;
		fir_coeff[117] = 16'hFF88;
		fir_coeff[118] = 16'hFF6A;
		fir_coeff[119] = 16'hFF8B;
		fir_coeff[120] = 16'hFFD6;
		fir_coeff[121] = 16'h2A;
		fir_coeff[122] = 16'h63;
		fir_coeff[123] = 16'h6F;
		fir_coeff[124] = 16'h4D;
		fir_coeff[125] = 16'h10;
		fir_coeff[126] = 16'hFFD2;
		fir_coeff[127] = 16'hFFAC;
		fir_coeff[128] = 16'hFFAC;
		fir_coeff[129] = 16'hFFCE;
		fir_coeff[130] = 16'h1;
		fir_coeff[131] = 16'h2F;
		fir_coeff[132] = 16'h46;
		fir_coeff[133] = 16'h3F;
		fir_coeff[134] = 16'h1F;
		fir_coeff[135] = 16'hFFF5;
		fir_coeff[136] = 16'hFFD3;
		fir_coeff[137] = 16'hFFC6;
		fir_coeff[138] = 16'hFFD1;
		fir_coeff[139] = 16'hFFEF;
		fir_coeff[140] = 16'h11;
		fir_coeff[141] = 16'h2A;
		fir_coeff[142] = 16'h30;
		fir_coeff[143] = 16'h22;
		fir_coeff[144] = 16'h7;
		fir_coeff[145] = 16'hFFEC;
		fir_coeff[146] = 16'hFFDB;
		fir_coeff[147] = 16'hFFDA;
		fir_coeff[148] = 16'hFFE9;
		fir_coeff[149] = 16'h0;
		fir_coeff[150] = 16'h15;
		fir_coeff[151] = 16'h20;
		fir_coeff[152] = 16'h1E;
		fir_coeff[153] = 16'hF;
		fir_coeff[154] = 16'hFFFC;
		fir_coeff[155] = 16'hFFEB;
		fir_coeff[156] = 16'hFFE5;
		fir_coeff[157] = 16'hFFE9;
		fir_coeff[158] = 16'hFFF7;
		fir_coeff[159] = 16'h7;
		fir_coeff[160] = 16'h13;
		fir_coeff[161] = 16'h17;
		fir_coeff[162] = 16'h11;
		fir_coeff[163] = 16'h5;
		fir_coeff[164] = 16'hFFF8;
		fir_coeff[165] = 16'hFFEF;
		fir_coeff[166] = 16'hFFEE;
		fir_coeff[167] = 16'hFFF4;
		fir_coeff[168] = 16'hFFFF;
		fir_coeff[169] = 16'h9;
		fir_coeff[170] = 16'hF;
		fir_coeff[171] = 16'hE;
		fir_coeff[172] = 16'h8;
		fir_coeff[173] = 16'hFFFF;
		fir_coeff[174] = 16'hFFF7;
		fir_coeff[175] = 16'hFFF3;
		fir_coeff[176] = 16'hFFF5;
		fir_coeff[177] = 16'hFFFB;
		fir_coeff[178] = 16'h2;
		fir_coeff[179] = 16'h8;
		fir_coeff[180] = 16'hB;
		fir_coeff[181] = 16'h9;
		fir_coeff[182] = 16'h3;
		fir_coeff[183] = 16'hFFFD;
		fir_coeff[184] = 16'hFFF8;
		fir_coeff[185] = 16'hFFF7;
		fir_coeff[186] = 16'hFFF9;
		fir_coeff[187] = 16'hFFFE;
		fir_coeff[188] = 16'h4;
		fir_coeff[189] = 16'h8;
		fir_coeff[190] = 16'h9;
		fir_coeff[191] = 16'h7;
		fir_coeff[192] = 16'h2;
		fir_coeff[193] = 16'hFFFC;
		fir_coeff[194] = 16'hFFF6;
		fir_coeff[195] = 16'hFFF2;
		fir_coeff[196] = 16'hFFF1;
		fir_coeff[197] = 16'hFFF2;
		fir_coeff[198] = 16'hFFF4;
		fir_coeff[199] = 16'hFFF8;
		fir_coeff[200] = 16'hFFFB;
		fir_coeff[201] = 16'hFFFE;
		fir_coeff[202] = 16'hFFFF;
		fir_coeff[203] = 16'h0;
	end
endmodule