// serves to load the coefficients for synthesis.
module coeff_broadcaster;
	reg  [15:0] fir_coeff [0:`FILTER_SIZE-1];

	initial begin
		fir_coeff[0] = 16'h1;
		fir_coeff[1] = 16'hFFFD;
		fir_coeff[2] = 16'hFFF7;
		fir_coeff[3] = 16'hFFED;
		fir_coeff[4] = 16'hFFE0;
		fir_coeff[5] = 16'hFFD2;
		fir_coeff[6] = 16'hFFC7;
		fir_coeff[7] = 16'hFFC3;
		fir_coeff[8] = 16'hFFC8;
		fir_coeff[9] = 16'hFFD8;
		fir_coeff[10] = 16'hFFEE;
		fir_coeff[11] = 16'h7;
		fir_coeff[12] = 16'h1B;
		fir_coeff[13] = 16'h24;
		fir_coeff[14] = 16'h20;
		fir_coeff[15] = 16'hF;
		fir_coeff[16] = 16'hFFF8;
		fir_coeff[17] = 16'hFFE5;
		fir_coeff[18] = 16'hFFDB;
		fir_coeff[19] = 16'hFFE1;
		fir_coeff[20] = 16'hFFF4;
		fir_coeff[21] = 16'hD;
		fir_coeff[22] = 16'h22;
		fir_coeff[23] = 16'h2A;
		fir_coeff[24] = 16'h21;
		fir_coeff[25] = 16'h8;
		fir_coeff[26] = 16'hFFEA;
		fir_coeff[27] = 16'hFFD3;
		fir_coeff[28] = 16'hFFCE;
		fir_coeff[29] = 16'hFFDD;
		fir_coeff[30] = 16'hFFFD;
		fir_coeff[31] = 16'h21;
		fir_coeff[32] = 16'h3A;
		fir_coeff[33] = 16'h3B;
		fir_coeff[34] = 16'h24;
		fir_coeff[35] = 16'hFFFA;
		fir_coeff[36] = 16'hFFD0;
		fir_coeff[37] = 16'hFFB7;
		fir_coeff[38] = 16'hFFBB;
		fir_coeff[39] = 16'hFFDE;
		fir_coeff[40] = 16'h13;
		fir_coeff[41] = 16'h43;
		fir_coeff[42] = 16'h5B;
		fir_coeff[43] = 16'h4D;
		fir_coeff[44] = 16'h1C;
		fir_coeff[45] = 16'hFFDB;
		fir_coeff[46] = 16'hFFA5;
		fir_coeff[47] = 16'hFF92;
		fir_coeff[48] = 16'hFFAE;
		fir_coeff[49] = 16'hFFEF;
		fir_coeff[50] = 16'h3E;
		fir_coeff[51] = 16'h77;
		fir_coeff[52] = 16'h82;
		fir_coeff[53] = 16'h54;
		fir_coeff[54] = 16'hFFFE;
		fir_coeff[55] = 16'hFFA2;
		fir_coeff[56] = 16'hFF67;
		fir_coeff[57] = 16'hFF6B;
		fir_coeff[58] = 16'hFFB0;
		fir_coeff[59] = 16'h1E;
		fir_coeff[60] = 16'h87;
		fir_coeff[61] = 16'hBF;
		fir_coeff[62] = 16'hA7;
		fir_coeff[63] = 16'h44;
		fir_coeff[64] = 16'hFFBB;
		fir_coeff[65] = 16'hFF45;
		fir_coeff[66] = 16'hFF17;
		fir_coeff[67] = 16'hFF4B;
		fir_coeff[68] = 16'hFFD4;
		fir_coeff[69] = 16'h7C;
		fir_coeff[70] = 16'hFD;
		fir_coeff[71] = 16'h119;
		fir_coeff[72] = 16'hBC;
		fir_coeff[73] = 16'h3;
		fir_coeff[74] = 16'hFF37;
		fir_coeff[75] = 16'hFEB0;
		fir_coeff[76] = 16'hFEB1;
		fir_coeff[77] = 16'hFF47;
		fir_coeff[78] = 16'h3E;
		fir_coeff[79] = 16'h135;
		fir_coeff[80] = 16'h1BD;
		fir_coeff[81] = 16'h18E;
		fir_coeff[82] = 16'hA7;
		fir_coeff[83] = 16'hFF59;
		fir_coeff[84] = 16'hFE2A;
		fir_coeff[85] = 16'hFDA7;
		fir_coeff[86] = 16'hFE22;
		fir_coeff[87] = 16'hFF88;
		fir_coeff[88] = 16'h15F;
		fir_coeff[89] = 16'h2E5;
		fir_coeff[90] = 16'h35C;
		fir_coeff[91] = 16'h25B;
		fir_coeff[92] = 16'h6;
		fir_coeff[93] = 16'hFD1D;
		fir_coeff[94] = 16'hFACB;
		fir_coeff[95] = 16'hFA4B;
		fir_coeff[96] = 16'hFC78;
		fir_coeff[97] = 16'h176;
		fir_coeff[98] = 16'h887;
		fir_coeff[99] = 16'h1039;
		fir_coeff[100] = 16'h16BF;
		fir_coeff[101] = 16'h1A7C;
		fir_coeff[102] = 16'h1A7C;
		fir_coeff[103] = 16'h16BF;
		fir_coeff[104] = 16'h1039;
		fir_coeff[105] = 16'h887;
		fir_coeff[106] = 16'h176;
		fir_coeff[107] = 16'hFC78;
		fir_coeff[108] = 16'hFA4B;
		fir_coeff[109] = 16'hFACB;
		fir_coeff[110] = 16'hFD1D;
		fir_coeff[111] = 16'h6;
		fir_coeff[112] = 16'h25B;
		fir_coeff[113] = 16'h35C;
		fir_coeff[114] = 16'h2E5;
		fir_coeff[115] = 16'h15F;
		fir_coeff[116] = 16'hFF88;
		fir_coeff[117] = 16'hFE22;
		fir_coeff[118] = 16'hFDA7;
		fir_coeff[119] = 16'hFE2A;
		fir_coeff[120] = 16'hFF59;
		fir_coeff[121] = 16'hA7;
		fir_coeff[122] = 16'h18E;
		fir_coeff[123] = 16'h1BD;
		fir_coeff[124] = 16'h135;
		fir_coeff[125] = 16'h3E;
		fir_coeff[126] = 16'hFF47;
		fir_coeff[127] = 16'hFEB1;
		fir_coeff[128] = 16'hFEB0;
		fir_coeff[129] = 16'hFF37;
		fir_coeff[130] = 16'h3;
		fir_coeff[131] = 16'hBC;
		fir_coeff[132] = 16'h119;
		fir_coeff[133] = 16'hFD;
		fir_coeff[134] = 16'h7C;
		fir_coeff[135] = 16'hFFD4;
		fir_coeff[136] = 16'hFF4B;
		fir_coeff[137] = 16'hFF17;
		fir_coeff[138] = 16'hFF45;
		fir_coeff[139] = 16'hFFBB;
		fir_coeff[140] = 16'h44;
		fir_coeff[141] = 16'hA7;
		fir_coeff[142] = 16'hBF;
		fir_coeff[143] = 16'h87;
		fir_coeff[144] = 16'h1E;
		fir_coeff[145] = 16'hFFB0;
		fir_coeff[146] = 16'hFF6B;
		fir_coeff[147] = 16'hFF67;
		fir_coeff[148] = 16'hFFA2;
		fir_coeff[149] = 16'hFFFE;
		fir_coeff[150] = 16'h54;
		fir_coeff[151] = 16'h82;
		fir_coeff[152] = 16'h77;
		fir_coeff[153] = 16'h3E;
		fir_coeff[154] = 16'hFFEF;
		fir_coeff[155] = 16'hFFAE;
		fir_coeff[156] = 16'hFF92;
		fir_coeff[157] = 16'hFFA5;
		fir_coeff[158] = 16'hFFDB;
		fir_coeff[159] = 16'h1C;
		fir_coeff[160] = 16'h4D;
		fir_coeff[161] = 16'h5B;
		fir_coeff[162] = 16'h43;
		fir_coeff[163] = 16'h13;
		fir_coeff[164] = 16'hFFDE;
		fir_coeff[165] = 16'hFFBB;
		fir_coeff[166] = 16'hFFB7;
		fir_coeff[167] = 16'hFFD0;
		fir_coeff[168] = 16'hFFFA;
		fir_coeff[169] = 16'h24;
		fir_coeff[170] = 16'h3B;
		fir_coeff[171] = 16'h3A;
		fir_coeff[172] = 16'h21;
		fir_coeff[173] = 16'hFFFD;
		fir_coeff[174] = 16'hFFDD;
		fir_coeff[175] = 16'hFFCE;
		fir_coeff[176] = 16'hFFD3;
		fir_coeff[177] = 16'hFFEA;
		fir_coeff[178] = 16'h8;
		fir_coeff[179] = 16'h21;
		fir_coeff[180] = 16'h2A;
		fir_coeff[181] = 16'h22;
		fir_coeff[182] = 16'hD;
		fir_coeff[183] = 16'hFFF4;
		fir_coeff[184] = 16'hFFE1;
		fir_coeff[185] = 16'hFFDB;
		fir_coeff[186] = 16'hFFE5;
		fir_coeff[187] = 16'hFFF8;
		fir_coeff[188] = 16'hF;
		fir_coeff[189] = 16'h20;
		fir_coeff[190] = 16'h24;
		fir_coeff[191] = 16'h1B;
		fir_coeff[192] = 16'h7;
		fir_coeff[193] = 16'hFFEE;
		fir_coeff[194] = 16'hFFD8;
		fir_coeff[195] = 16'hFFC8;
		fir_coeff[196] = 16'hFFC3;
		fir_coeff[197] = 16'hFFC7;
		fir_coeff[198] = 16'hFFD2;
		fir_coeff[199] = 16'hFFE0;
		fir_coeff[200] = 16'hFFED;
		fir_coeff[201] = 16'hFFF7;
		fir_coeff[202] = 16'hFFFD;
		fir_coeff[203] = 16'h1;
	end
endmodule