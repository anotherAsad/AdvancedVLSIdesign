power['h0] = 'h1;		log['h0] = 'hf;
power['h1] = 'h2;		log['h1] = 'h0;
power['h2] = 'h4;		log['h2] = 'h1;
power['h3] = 'h8;		log['h3] = 'h19;
power['h4] = 'h10;		log['h4] = 'h2;
power['h5] = 'h20;		log['h5] = 'h32;
power['h6] = 'h40;		log['h6] = 'h1a;
power['h7] = 'h80;		log['h7] = 'hc6;
power['h8] = 'h1d;		log['h8] = 'h3;
power['h9] = 'h3a;		log['h9] = 'hdf;
power['ha] = 'h74;		log['ha] = 'h33;
power['hb] = 'he8;		log['hb] = 'hee;
power['hc] = 'hcd;		log['hc] = 'h1b;
power['hd] = 'h87;		log['hd] = 'h68;
power['he] = 'h13;		log['he] = 'hc7;
power['hf] = 'h26;		log['hf] = 'h4b;
power['h10] = 'h4c;		log['h10] = 'h4;
power['h11] = 'h98;		log['h11] = 'h64;
power['h12] = 'h2d;		log['h12] = 'he0;
power['h13] = 'h5a;		log['h13] = 'he;
power['h14] = 'hb4;		log['h14] = 'h34;
power['h15] = 'h75;		log['h15] = 'h8d;
power['h16] = 'hea;		log['h16] = 'hef;
power['h17] = 'hc9;		log['h17] = 'h81;
power['h18] = 'h8f;		log['h18] = 'h1c;
power['h19] = 'h3;		log['h19] = 'hc1;
power['h1a] = 'h6;		log['h1a] = 'h69;
power['h1b] = 'hc;		log['h1b] = 'hf8;
power['h1c] = 'h18;		log['h1c] = 'hc8;
power['h1d] = 'h30;		log['h1d] = 'h8;
power['h1e] = 'h60;		log['h1e] = 'h4c;
power['h1f] = 'hc0;		log['h1f] = 'h71;
power['h20] = 'h9d;		log['h20] = 'h5;
power['h21] = 'h27;		log['h21] = 'h8a;
power['h22] = 'h4e;		log['h22] = 'h65;
power['h23] = 'h9c;		log['h23] = 'h2f;
power['h24] = 'h25;		log['h24] = 'he1;
power['h25] = 'h4a;		log['h25] = 'h24;
power['h26] = 'h94;		log['h26] = 'hf;
power['h27] = 'h35;		log['h27] = 'h21;
power['h28] = 'h6a;		log['h28] = 'h35;
power['h29] = 'hd4;		log['h29] = 'h93;
power['h2a] = 'hb5;		log['h2a] = 'h8e;
power['h2b] = 'h77;		log['h2b] = 'hda;
power['h2c] = 'hee;		log['h2c] = 'hf0;
power['h2d] = 'hc1;		log['h2d] = 'h12;
power['h2e] = 'h9f;		log['h2e] = 'h82;
power['h2f] = 'h23;		log['h2f] = 'h45;
power['h30] = 'h46;		log['h30] = 'h1d;
power['h31] = 'h8c;		log['h31] = 'hb5;
power['h32] = 'h5;		log['h32] = 'hc2;
power['h33] = 'ha;		log['h33] = 'h7d;
power['h34] = 'h14;		log['h34] = 'h6a;
power['h35] = 'h28;		log['h35] = 'h27;
power['h36] = 'h50;		log['h36] = 'hf9;
power['h37] = 'ha0;		log['h37] = 'hb9;
power['h38] = 'h5d;		log['h38] = 'hc9;
power['h39] = 'hba;		log['h39] = 'h9a;
power['h3a] = 'h69;		log['h3a] = 'h9;
power['h3b] = 'hd2;		log['h3b] = 'h78;
power['h3c] = 'hb9;		log['h3c] = 'h4d;
power['h3d] = 'h6f;		log['h3d] = 'he4;
power['h3e] = 'hde;		log['h3e] = 'h72;
power['h3f] = 'ha1;		log['h3f] = 'ha6;
power['h40] = 'h5f;		log['h40] = 'h6;
power['h41] = 'hbe;		log['h41] = 'hbf;
power['h42] = 'h61;		log['h42] = 'h8b;
power['h43] = 'hc2;		log['h43] = 'h62;
power['h44] = 'h99;		log['h44] = 'h66;
power['h45] = 'h2f;		log['h45] = 'hdd;
power['h46] = 'h5e;		log['h46] = 'h30;
power['h47] = 'hbc;		log['h47] = 'hfd;
power['h48] = 'h65;		log['h48] = 'he2;
power['h49] = 'hca;		log['h49] = 'h98;
power['h4a] = 'h89;		log['h4a] = 'h25;
power['h4b] = 'hf;		log['h4b] = 'hb3;
power['h4c] = 'h1e;		log['h4c] = 'h10;
power['h4d] = 'h3c;		log['h4d] = 'h91;
power['h4e] = 'h78;		log['h4e] = 'h22;
power['h4f] = 'hf0;		log['h4f] = 'h88;
power['h50] = 'hfd;		log['h50] = 'h36;
power['h51] = 'he7;		log['h51] = 'hd0;
power['h52] = 'hd3;		log['h52] = 'h94;
power['h53] = 'hbb;		log['h53] = 'hce;
power['h54] = 'h6b;		log['h54] = 'h8f;
power['h55] = 'hd6;		log['h55] = 'h96;
power['h56] = 'hb1;		log['h56] = 'hdb;
power['h57] = 'h7f;		log['h57] = 'hbd;
power['h58] = 'hfe;		log['h58] = 'hf1;
power['h59] = 'he1;		log['h59] = 'hd2;
power['h5a] = 'hdf;		log['h5a] = 'h13;
power['h5b] = 'ha3;		log['h5b] = 'h5c;
power['h5c] = 'h5b;		log['h5c] = 'h83;
power['h5d] = 'hb6;		log['h5d] = 'h38;
power['h5e] = 'h71;		log['h5e] = 'h46;
power['h5f] = 'he2;		log['h5f] = 'h40;
power['h60] = 'hd9;		log['h60] = 'h1e;
power['h61] = 'haf;		log['h61] = 'h42;
power['h62] = 'h43;		log['h62] = 'hb6;
power['h63] = 'h86;		log['h63] = 'ha3;
power['h64] = 'h11;		log['h64] = 'hc3;
power['h65] = 'h22;		log['h65] = 'h48;
power['h66] = 'h44;		log['h66] = 'h7e;
power['h67] = 'h88;		log['h67] = 'h6e;
power['h68] = 'hd;		log['h68] = 'h6b;
power['h69] = 'h1a;		log['h69] = 'h3a;
power['h6a] = 'h34;		log['h6a] = 'h28;
power['h6b] = 'h68;		log['h6b] = 'h54;
power['h6c] = 'hd0;		log['h6c] = 'hfa;
power['h6d] = 'hbd;		log['h6d] = 'h85;
power['h6e] = 'h67;		log['h6e] = 'hba;
power['h6f] = 'hce;		log['h6f] = 'h3d;
power['h70] = 'h81;		log['h70] = 'hca;
power['h71] = 'h1f;		log['h71] = 'h5e;
power['h72] = 'h3e;		log['h72] = 'h9b;
power['h73] = 'h7c;		log['h73] = 'h9f;
power['h74] = 'hf8;		log['h74] = 'ha;
power['h75] = 'hed;		log['h75] = 'h15;
power['h76] = 'hc7;		log['h76] = 'h79;
power['h77] = 'h93;		log['h77] = 'h2b;
power['h78] = 'h3b;		log['h78] = 'h4e;
power['h79] = 'h76;		log['h79] = 'hd4;
power['h7a] = 'hec;		log['h7a] = 'he5;
power['h7b] = 'hc5;		log['h7b] = 'hac;
power['h7c] = 'h97;		log['h7c] = 'h73;
power['h7d] = 'h33;		log['h7d] = 'hf3;
power['h7e] = 'h66;		log['h7e] = 'ha7;
power['h7f] = 'hcc;		log['h7f] = 'h57;
power['h80] = 'h85;		log['h80] = 'h7;
power['h81] = 'h17;		log['h81] = 'h70;
power['h82] = 'h2e;		log['h82] = 'hc0;
power['h83] = 'h5c;		log['h83] = 'hf7;
power['h84] = 'hb8;		log['h84] = 'h8c;
power['h85] = 'h6d;		log['h85] = 'h80;
power['h86] = 'hda;		log['h86] = 'h63;
power['h87] = 'ha9;		log['h87] = 'hd;
power['h88] = 'h4f;		log['h88] = 'h67;
power['h89] = 'h9e;		log['h89] = 'h4a;
power['h8a] = 'h21;		log['h8a] = 'hde;
power['h8b] = 'h42;		log['h8b] = 'hed;
power['h8c] = 'h84;		log['h8c] = 'h31;
power['h8d] = 'h15;		log['h8d] = 'hc5;
power['h8e] = 'h2a;		log['h8e] = 'hfe;
power['h8f] = 'h54;		log['h8f] = 'h18;
power['h90] = 'ha8;		log['h90] = 'he3;
power['h91] = 'h4d;		log['h91] = 'ha5;
power['h92] = 'h9a;		log['h92] = 'h99;
power['h93] = 'h29;		log['h93] = 'h77;
power['h94] = 'h52;		log['h94] = 'h26;
power['h95] = 'ha4;		log['h95] = 'hb8;
power['h96] = 'h55;		log['h96] = 'hb4;
power['h97] = 'haa;		log['h97] = 'h7c;
power['h98] = 'h49;		log['h98] = 'h11;
power['h99] = 'h92;		log['h99] = 'h44;
power['h9a] = 'h39;		log['h9a] = 'h92;
power['h9b] = 'h72;		log['h9b] = 'hd9;
power['h9c] = 'he4;		log['h9c] = 'h23;
power['h9d] = 'hd5;		log['h9d] = 'h20;
power['h9e] = 'hb7;		log['h9e] = 'h89;
power['h9f] = 'h73;		log['h9f] = 'h2e;
power['ha0] = 'he6;		log['ha0] = 'h37;
power['ha1] = 'hd1;		log['ha1] = 'h3f;
power['ha2] = 'hbf;		log['ha2] = 'hd1;
power['ha3] = 'h63;		log['ha3] = 'h5b;
power['ha4] = 'hc6;		log['ha4] = 'h95;
power['ha5] = 'h91;		log['ha5] = 'hbc;
power['ha6] = 'h3f;		log['ha6] = 'hcf;
power['ha7] = 'h7e;		log['ha7] = 'hcd;
power['ha8] = 'hfc;		log['ha8] = 'h90;
power['ha9] = 'he5;		log['ha9] = 'h87;
power['haa] = 'hd7;		log['haa] = 'h97;
power['hab] = 'hb3;		log['hab] = 'hb2;
power['hac] = 'h7b;		log['hac] = 'hdc;
power['had] = 'hf6;		log['had] = 'hfc;
power['hae] = 'hf1;		log['hae] = 'hbe;
power['haf] = 'hff;		log['haf] = 'h61;
power['hb0] = 'he3;		log['hb0] = 'hf2;
power['hb1] = 'hdb;		log['hb1] = 'h56;
power['hb2] = 'hab;		log['hb2] = 'hd3;
power['hb3] = 'h4b;		log['hb3] = 'hab;
power['hb4] = 'h96;		log['hb4] = 'h14;
power['hb5] = 'h31;		log['hb5] = 'h2a;
power['hb6] = 'h62;		log['hb6] = 'h5d;
power['hb7] = 'hc4;		log['hb7] = 'h9e;
power['hb8] = 'h95;		log['hb8] = 'h84;
power['hb9] = 'h37;		log['hb9] = 'h3c;
power['hba] = 'h6e;		log['hba] = 'h39;
power['hbb] = 'hdc;		log['hbb] = 'h53;
power['hbc] = 'ha5;		log['hbc] = 'h47;
power['hbd] = 'h57;		log['hbd] = 'h6d;
power['hbe] = 'hae;		log['hbe] = 'h41;
power['hbf] = 'h41;		log['hbf] = 'ha2;
power['hc0] = 'h82;		log['hc0] = 'h1f;
power['hc1] = 'h19;		log['hc1] = 'h2d;
power['hc2] = 'h32;		log['hc2] = 'h43;
power['hc3] = 'h64;		log['hc3] = 'hd8;
power['hc4] = 'hc8;		log['hc4] = 'hb7;
power['hc5] = 'h8d;		log['hc5] = 'h7b;
power['hc6] = 'h7;		log['hc6] = 'ha4;
power['hc7] = 'he;		log['hc7] = 'h76;
power['hc8] = 'h1c;		log['hc8] = 'hc4;
power['hc9] = 'h38;		log['hc9] = 'h17;
power['hca] = 'h70;		log['hca] = 'h49;
power['hcb] = 'he0;		log['hcb] = 'hec;
power['hcc] = 'hdd;		log['hcc] = 'h7f;
power['hcd] = 'ha7;		log['hcd] = 'hc;
power['hce] = 'h53;		log['hce] = 'h6f;
power['hcf] = 'ha6;		log['hcf] = 'hf6;
power['hd0] = 'h51;		log['hd0] = 'h6c;
power['hd1] = 'ha2;		log['hd1] = 'ha1;
power['hd2] = 'h59;		log['hd2] = 'h3b;
power['hd3] = 'hb2;		log['hd3] = 'h52;
power['hd4] = 'h79;		log['hd4] = 'h29;
power['hd5] = 'hf2;		log['hd5] = 'h9d;
power['hd6] = 'hf9;		log['hd6] = 'h55;
power['hd7] = 'hef;		log['hd7] = 'haa;
power['hd8] = 'hc3;		log['hd8] = 'hfb;
power['hd9] = 'h9b;		log['hd9] = 'h60;
power['hda] = 'h2b;		log['hda] = 'h86;
power['hdb] = 'h56;		log['hdb] = 'hb1;
power['hdc] = 'hac;		log['hdc] = 'hbb;
power['hdd] = 'h45;		log['hdd] = 'hcc;
power['hde] = 'h8a;		log['hde] = 'h3e;
power['hdf] = 'h9;		log['hdf] = 'h5a;
power['he0] = 'h12;		log['he0] = 'hcb;
power['he1] = 'h24;		log['he1] = 'h59;
power['he2] = 'h48;		log['he2] = 'h5f;
power['he3] = 'h90;		log['he3] = 'hb0;
power['he4] = 'h3d;		log['he4] = 'h9c;
power['he5] = 'h7a;		log['he5] = 'ha9;
power['he6] = 'hf4;		log['he6] = 'ha0;
power['he7] = 'hf5;		log['he7] = 'h51;
power['he8] = 'hf7;		log['he8] = 'hb;
power['he9] = 'hf3;		log['he9] = 'hf5;
power['hea] = 'hfb;		log['hea] = 'h16;
power['heb] = 'heb;		log['heb] = 'heb;
power['hec] = 'hcb;		log['hec] = 'h7a;
power['hed] = 'h8b;		log['hed] = 'h75;
power['hee] = 'hb;		log['hee] = 'h2c;
power['hef] = 'h16;		log['hef] = 'hd7;
power['hf0] = 'h2c;		log['hf0] = 'h4f;
power['hf1] = 'h58;		log['hf1] = 'hae;
power['hf2] = 'hb0;		log['hf2] = 'hd5;
power['hf3] = 'h7d;		log['hf3] = 'he9;
power['hf4] = 'hfa;		log['hf4] = 'he6;
power['hf5] = 'he9;		log['hf5] = 'he7;
power['hf6] = 'hcf;		log['hf6] = 'had;
power['hf7] = 'h83;		log['hf7] = 'he8;
power['hf8] = 'h1b;		log['hf8] = 'h74;
power['hf9] = 'h36;		log['hf9] = 'hd6;
power['hfa] = 'h6c;		log['hfa] = 'hf4;
power['hfb] = 'hd8;		log['hfb] = 'hea;
power['hfc] = 'had;		log['hfc] = 'ha8;
power['hfd] = 'h47;		log['hfd] = 'h50;
power['hfe] = 'h8e;		log['hfe] = 'h58;
power['hff] = 'h1;		log['hff] = 'haf;